-- ****************************************
-- tittle:	Controlador para el ADS1115
-- author:	
-- date:		
-- description:
-- ****************************************